module cong(a,b);

input a;
output b;

assign a=~b;

endmodule;